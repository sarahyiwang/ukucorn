// Enabled counter with synchronous reset
module counter_en #(parameter N = 8)
					(input logic clk, reset, en,
					 output logic [N-1:0] q);
	always_ff@(posedge clk)
		if (reset)	q <= 0;
		else if (en) q <= q + 1;
endmodule

// Counter with async reset (non-enabled)
module counter #(parameter N = 8)
					(input logic clk, reset,
					 output logic [N-1:0] q);
	always_ff@(posedge clk, posedge reset)
		if (reset)	q <= 0;
		else q <= q + 1;
endmodule

/*
 * Address Generation Unit
 * Functions:
 *   1) Generate addresses for reading and writing of data RAM
 *   2) Retrieve twiddle factors
 *   3) Generate write signals for the data RAM
 * Keep track of:
 *   1) Which butterfly we are executing
 *   2) Which FFT level we are working on
 */ 

module AGU
	#(parameter logN = 9)
	(input logic clk, reset,
	 input logic StartFFT,
	 output logic FFTDone,
	 output logic [logN-1:0] MemA_Addr, MemB_Addr,
	 output logic [logN-2:0] TwAddr);
	
	logic [3:0] i; // Level of FFT counter
	logic [logN-2:0] j; // Butterfly index counter
	logic [logN-1:0] ja, jb; // For calculating addresses
	logic [1:0] k; // Wait until A' and B' are written to memory

	// Synchronize StartFFT and assert ClearHold
	logic StartFFT1;
	logic ClearHold;
	
	always_ff @(posedge clk)
			StartFFT1 <= StartFFT;
			
	assign ClearHold = StartFFT & ~StartFFT1;

	counter_en #(4) fft_counter(clk, i_reset, i_en, i); // FFT Level counter
	counter_en #(logN-1) butterfly_counter(clk, j_reset, j_en, j); // Butterfly index counter
	counter_en #(2) hold_counter(clk, k_reset, k_en, k); // Hold counter
	
	assign i_reset = ClearHold | (i == logN); // reset when maxed out
	assign j_reset = ClearHold | (&k); // reset when k is maxed out
	assign k_reset = ClearHold | &k; // reset when maxed out
	
	assign i_en = &k; // enable when k is maxed out
	assign j_en = ~(&j); // enable while not maxed out
	assign k_en = &j; // enable when j is maxed out
	
	// Generate addresses for data and twiddles
	assign ja = j << 1;
	assign jb = ja + 1;
	assign MemA_Addr = (ja << i) | (ja >> (logN - i));
	assign MemB_Addr = (jb << i) | (jb >> (logN - i));
	
	// Twiddle mask generator - a right shift register
	// that fills up with 1s as the level counter is incremented
	logic [logN-2:0] ones = ~0;
	logic [logN-2:0] zeros = 0;
	assign TwAddr = ({ones, zeros} >> i) & j;
	
	always_ff @(posedge clk) begin
	  if (ClearHold) FFTDone <= 0;
	  else if (&k & (i == logN)) FFTDone <= 1;
	end
endmodule // agu

/*
 * http://www.cs.columbia.edu/~sedwards/classes/2015/4840/memory.pdf
 */
module TwoPortRAM
	#(parameter logN)
	(input logic clk,
	 input logic [logN-1:0] AddA, AddB, // address
	 input logic [31:0] Ain, Bin, // data in
	 input logic WriteA, WriteB, // write enables
	 output logic [31:0] Aout, Bout);

	parameter N = 1 << logN;
	logic [31:0] Mem [N-1:0];

	always_ff @(posedge clk) begin
		if (WriteA) begin
			Mem[AddA] <= Ain;
			Aout <= Ain; end
		else Aout <= Mem[AddA]; end

	always_ff @(posedge clk) begin
		if (WriteB) begin
			Mem[AddB] <= Bin;
			Bout <= Bin; end
		else Bout <= Mem[AddB]; end
endmodule // TwoPortRAM


module BFU
	#(parameter logN = 9)
	(input logic [15:0] A_r, A_i, // A
	 input logic [15:0] B_r, B_i, // B
	 input logic signed [15:0] Tw_r, Tw_i, // Tw_r = TwV_real[TwAddr]
	 output logic signed [15:0] Ap_r, Ap_i,  // A'
	 output logic signed [15:0] Bp_r, Bp_i); // B'

	logic signed [31:0] temp_r, temp_i;
	logic signed [15:0] temp_r_p, temp_i_p; // pruned version of T1

	// Complex multiplier
	assign temp_r = (B_r * Tw_r) - (B_i * Tw_i);
	assign temp_i = (B_r * Tw_i) + (B_i * Tw_r);

	// Prune T1
	assign temp_r_p = temp_r[30:15];
	assign temp_i_p = temp_i[30:15];

	// Complex adder for A'
	assign Ap_r = A_r + temp_r_p;
	assign Ap_i = A_i + temp_i_p;

	// Complex adder for B'
	assign Bp_r = A_r - temp_r_p;
	assign Bp_i = A_i - temp_i_p;
endmodule // BFU

module ukucorn
	#(parameter logN = 9)
	(input logic clk, reset,
	 input logic [10:0] data);

	//////////////////////////////////////
	//////          STATES          //////
	//////////////////////////////////////
	
	// idle: nothing to do...
	// sample: take data from ADC
	// load: load samples into RAM
	// fft: process data
	// find_freq: find the four dominant frequencies
	logic [2:0] state, nextstate;
	typedef enum logic [2:0] {idle, sample, load, fft, find} statetype;
	
	// Next state register
	always_ff @(posedge clk, posedge reset)
		begin
			if (reset) state <= idle;
			else state <= nextstate;
		end
	 
	//////////////////////////////////////
	//////       SAMPLE DATA        //////
	//////////////////////////////////////
	
	parameter threshold = 0;
	logic [logN-1:0] sample_count;
	logic sc_reset;
	assign sc_reset = ~(state == sample); // suppress counter when not in sample state
	counter #(logN) sample_counter(clk, sc_reset, sample_count);

	//////////////////////////////////////
	//////        LOAD DATA         //////
	//////////////////////////////////////

	logic LoadWrite;
	assign LoadWrite = (state == load); // enable write to memory
	logic [logN-2:0] load_count;
	logic lc_reset;
	assign lc_reset = ~LoadWrite; // suppress counter when not in sample stat
	counter #(logN-1) load_counter(clk, lc_reset, load_count);

	logic [logN-1:0] a0, a1; // write 2 data points at once
	
	// Load address counter
	always_ff @(posedge clk, posedge reset)
		if (reset) begin
			a0 <= 0; a1 <= 1; end
		else if (LoadWrite) begin
			a0 <= a0 + 2;
			a1 <= a1 + 2; end

	//////////////////////////////////////
	//////            FFT           ////// 
	//////////////////////////////////////

	// AGU signals
	logic StartFFT, FFTDone;
	logic FFTWrite, MemWrite;
	logic [logN-1:0] ja, jb;
	logic [logN-2:0] TwAddr;

	// BFU signals
	logic signed [15:0] Tw_r, Tw_i;
	logic signed [15:0] A_r, A_i;
	logic signed [15:0] B_r, B_i;
	logic signed [15:0] Ap_r, Ap_i;
	logic signed [15:0] Bp_r, Bp_i;

	// RAM signals
	logic [logN-1:0] MemA_Addr, MemB_Addr;
	logic [31:0] Ain, Aout, Bin, Bout;

	// Divide the clock by 2 (read, write)
	logic rwclk;
	logic [1:0] q;
	counter #(2) clk_counter(clk, reset, q);
	assign rwclk = q[1]; // read: 10; write: 11
	assign FFTRead = (q == 2'b11) & (state == fft);
	assign FFTWrite = (q == 2'b00) & (state == fft);
	assign StartFFT = (state == fft);
 	
	AGU #(logN) agu1(rwclk, reset, StartFFT, FFTDone, ja, jb, TwAddr);
	BFU #(logN) bfu1(A_r, A_i, B_r, B_i, Tw_r, Tw_i, Ap_r, Ap_i, Bp_r, Bp_i);

	// To prevent timing errors, load A and B of BFU
	// only when FFTRead is high
	always_ff @(posedge FFTRead, posedge reset)
	 if (reset) begin
	    A_r <= 0;
		  A_i <= 0;
		  B_r <= 0;
		  B_i <= 0; end
	 else begin
		  A_r <= Aout[31:16];
		  A_i <= Aout[15:0];
		  B_r <= Bout[31:16];
		  B_i <= Bout[15:0];
	 end
	 
	logic [31:0] Ap, Bp;
	
	always_ff @(posedge FFTWrite, posedge reset)
	 if (reset) begin
	    Ap <= 0;
		  Bp <= 0; end
	 else begin
		  Ap <= {Ap_r, Ap_i};
		  Bp <= {Bp_r, Bp_i};
	 end
	
	
	assign MemWrite = FFTWrite | LoadWrite;
	assign MemA_Addr = LoadWrite ? a0 : ja;
	assign MemB_Addr = LoadWrite ? a1 : jb;

	TwoPortRAM #(logN) ram1(clk, MemA_Addr, MemB_Addr, Ain, Bin, MemWrite, MemWrite, Aout, Bout);

	// Twiddle Factor ROM
 	// Contains the look-up table of real and imaginary values
 	// of the required "roots of unity" that are passed to the BFU
 	parameter RomDepth = 1 << (logN -1); // N/2
 	logic [15:0] TwRom_r[0:RomDepth-1]; // 16-bit entries, N total
 	logic [15:0] TwRom_i[0:RomDepth-1];
 	initial $readmemh("Tw_r.txt",TwRom_r);
 	initial $readmemh("Tw_i.txt",TwRom_i);
 	
 	// Extract real and imaginary components
 	logic [15:0] zeros = 0;
	assign Tw_r = TwRom_r[TwAddr];
 	assign Tw_i = TwRom_i[TwAddr];
	assign Ain = LoadWrite ? {data, zeros} : Ap; // A'
	assign Bin = LoadWrite ? {zeros, zeros} : Bp;
	
	logic FindDone = 0;
	// Next state logic
	always_comb
	 case(state)
	    idle:	if (data > threshold) nextstate <= sample; // something detected!
	            else nextstate <= idle;
	    sample: if (&sample_count) nextstate <= load; // N samples reached
	            else nextstate <= sample;
	    load:   if (&load_count) nextstate <= fft; // 2 writes per cycle, so count up to N/2
	            else nextstate <= load;
	    fft:    if (FFTDone) nextstate <= find;
	            else nextstate <= fft;
	    find:   if (FindDone) nextstate <= find;
	            else nextstate <= fft;
	    default: nextstate <= idle;
	 endcase
 endmodule // main